module uart_tx ( 
);
endmodule