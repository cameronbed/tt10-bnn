// controller.v
// Handles state changes and control signals for the BNN
